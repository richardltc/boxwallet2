module app

// App
const app_name = 'BoxWallet Manager'
const app_version = '0.0.1'

pub fn name() string {
	return app_name
}

pub fn version() string {
	return app_version
}
